PK   �qU*4�
  �i     cirkitFile.json͜�n�8�_��a�Y9$�'߶w\��6�.��@�%�Α|�ܴ��e�ے,���I$�M�h4��pH�~�j�M�IZ�*���eQ���V�ٽ��L�EQ&M�|���ֻx0����B�iu��JU6I�i���g��|�8��Y&����*R3����fr�8ŉN��Ĺ?$���\0�GTJ��~���x���d�v��se�\9��,ĉG8�	+v$��;E�N9R^ ���pd��LIƴ`����B(?�b��N��H�9�,E�K��]�&j$��FB���L1?`$���ԟ�4�9�E*f�d�Գ��H�I= �d΅3��\���!�g��[��=gY] �L1W�G\0�#W��Ј+��q�1�ғ��8��FL��Ce����:$��U�\�x!��(�D8�h�FK�#�'�N��N�DN��n�s�z�|�~)w�����4t2*�������(���Pn(7���M&�h=�p��qC1sC1{�b���<a�8�`ۺ�������ȶ�>n�m��@˾-��v��Fa�R��ZΑ-^8�h�N�'Z'ZB'Z"'Zb7�9���������������������bp���Pn(7������bpC1������=K�uA���Ɩg�uA����Y�x-��肶Tߛ��lRd߽�h���Z&��LU��z��3U{W�7;��]T���kY̓,��1�2
�ϩ��T�ꀓ\�TeA���J���.�~��z7�[�LYTˮ)��#�C�F������}�,�G|v�FY�,!H�P+�_�)ǐ>9u�&V�:��(��Z�lV�:�W�5�,8�X,,�.�PG�8�f0�3G������"7�1��8���8�hr?9��9oc�l���S�W��ꛮ�d�*����o��1֠,r]>Yt��7[?:1�g��Gx�jo�뢲����� ��[���ּ/�(~Bi|��ש���U
e7�A�������LJN�������L�{��Q^d���3�3�x����tQ�*Y�p�2������~�bm��ohv����:�3�E�W�.�a�V��U��;.�1y���������N(n&��W�����>���۞�[��]�<o���<Cʛc���<f�ӆA!@�]�����1�.4�X>)P�%�=?�R �
����z�"��C��`:qb�l���}XN�)`9l�lO��|`�a9eXN�N���M��'��l}$�n��>g���ٍP��r#��>'70�q����)I����Im 3��6<��{c�׬+�*�6Կƅ���v4=��JM_j:Sӛ�����F�	0��6`$�]40�"�	0�H���6 u�75�E\wBZ���{�ݫ��K�''����+,�G��c �54ȳ*���+�I�a�A}y�p�p4�����p��ݨh��ݹ����Q����wf�m��a�4�a�4�al��)��do�(�*����;
r"�s#�� L�(J��#aD�$����Q���ǒ���CH!��y��CMXR�"�GA��L�=IJH��ZhY�=:F�W2���'�4��K1O���mc��כ��b�7٘��оtYWU7�j'��Ei���M]�f���w�i�x��|e����DtU�"�~����?��z��\ΗJ7.U��X��ھV���Ze�E��Q��N��\�ͪV�1���Y�ޞq`��Te�,����|E�P�Q7L���1����3[6�0?��!'�/	��h��+�97���Y�k��y�Uu��%��x-<iQ�s�	��$��}��I�<my��m	Gek�2lT��ʐ1�p�A���cГ���0��Q�u�#B'����]]�i����|j!t��Fc24��2|TFe�aڴD�hl���4�i���3��m-i�ϼ~ӎ���f�՗�o&��N�稱y�F�[ȁ���UѼ�Pf+#����!�bj<N����I@����:$t?5r�Ӏ��WQ>�l�+"u"3�E���V���hU��S�z��gG�4B���!�>���A&��X�1�#�_�!��Ӂ��??^�,�`���d�o�'̭�L#F`;fa�M!�݌��A2�Q?5�2�(�r?ω�t	@�L��d�(��i���.ᄱ���;m�Y��������He��xu��N�8!� ������J����ů�$�ަ:��&��������[�Ϊ�rgϮ�����8tٮ��оD�t��}�>�g���bJ�t��mu7S��O����̖G���ݳ�c$��lau�>�}4������A��"�gR2�p�BHa��9S�ed��
��x�����J�i�9��*�Z=E�Z�"Y��Q������ӹ}��3������x=�1y�Z�u�tRփ����/����l���Ve�ˠ�Z5͏/����|����p�2��.�����ڛ\�(��(?dm��;1�6UfGu����jy�٩mZ��ݙ�������m������3��O��i���4K��ŕ��-�]��f:L��,'����;u'�m���/��y��5r}|�v;|�ݬ�܅����,�9żS��F������Md�n�řu�����t�\���������#&�/l�I�7�d��^��ٴ;�G���#�������ǧ�M��>6������i��>v�5X�c�փ=>'�f��	�!�NMo+N�o�V�N1��i��m,@pN��"¬����S�Q6�.�T�r41��I��}��J��Wwu�47u��=�PK
   �qU*4�
  �i                   cirkitFile.jsonPK      =       