PK   LvU;��  �*     cirkitFile.json͚�r�6�_%C'w�����wuۙf�$�$�^x=�@"f�a�O������zĮ��]6J�N|�H::��ΏX�;����8�j�u�W�sF��\�Z��ݧ�u�y�U����k���ܣ�n�QZ�,�R�m�B�G�W(Lx�X�("4A�L�O0"?��svyl0fa���� :@�dP��
}I��?��{l,���"Q�a���3��a�0N��0,a⫣���&S��Y�4����5Q���(�Cɣ$Ȓ���Z3�2�5��l�a�g�4Մ���l�af�S�<F��c|��'�6���	KiUT�İ��i�C}<�؆	�,���Rl]�H�~#���}AJڌ�b늧Wd�V3�B?g#[�g�Bvl�Űie��bXꮭe1ÓR�1�.峺Xc8]�<���I��p������Ԯba��O�s�ۼ�M�,��U�4D��)��2����?�D5%�O�ndfKO����-wlR�}��^�o�� �,�1/A�o㕙|��<��S�yR�� ��O�A��]^n2���2g�޻\MM�x�odדּ�@�Ԫs ͟���F\ź �[�u%0�v�ڲֵ���,�7��VL�� �1|��gNn� �����6���:��Y��,��n��R�fY14���Mz�3�:���/Ǟ"�,d�mƓ[��Oz�6)�m)lMm^�D�C
�W�}f�p�D�D�躉6����eQ�I��J*�kP}eU\�Mk���Dc��&�EBP�}�S��L����;_~\謅#��%Y*S~���eYJ�O�x��q$�1�ݿ�F<��b#�]���g����]��R�m���u�,͗���i�� ���ܛV��(���Q����fpહ�n_�?�P�,�E�������ɓBo�����Y� ZX��,�L�mW����ݶj���6�*��C��m����Lx~�CFy�B�\F�'X���;��F� �ъdI�J��|���E(Y�I�~��r�ZY��1V9�u�:�ɕj���i��ƼDD���)����a��P�h��@�a��۶Sy���w	�x�À�1(��&_i�cUuf'7��鴱�xc���������\���~�]P\�(��	����0�*t=�V�m��g�k�
nvri6���G�G�#�������cu���:B�ȯ��D��^g���֜�o�wG�=%����j��� H��K�����(��G�A��\r���1&�0�rH�U�bE+���o��%��\s�U�~I #a�į���.o��(Ug��f�PF�� �"�]p����.��4`��!�iD9����F�TD��p��U):D��?\�G�&zE�e=(a�qy`����t0֑�����4������{ȉ�u%,g��H�á�u��F��Dz��)�%(�J�D1&3!��0��됨4�	�:�	Z�PC�D��2XX�t��w�?ˈ����1�WKS���`�{U��I�A��·�j��~0�������=�08
<���ħ�Ȼ=��)�k��7�E����}�o�0�MB�_8�K�s�x��i��F��E^�P}�W�za�T'Eٝ�zQ��};�j ���[Vy�^����u�X,SO��.L�������|�ak�U�k'J��^{5�N/!Nw�zX8�ɾ�W���is:����6�����WY�+�&�S6������'��dؽ��&d|�jߘ��LF	�~E���X�K��a�X�a�k�Al���&�rܚt���^#����bNO�јs{��Ɯ�����o��Ϻ�ø1��Y�x�����s��^��&�[��p���yu��7�Y�Ճ��PK
   LvU;��  �*                   cirkitFile.jsonPK      =   L    